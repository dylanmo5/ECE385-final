module top_pdm (
  input logic Clk,
  input logic reset_rtl_0,
  // TODO 
)
